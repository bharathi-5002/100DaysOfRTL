module excess_three_codes(x,y);
input [3:0]x;
output [3:0]y;
assign y = x + 3;
endmodule
